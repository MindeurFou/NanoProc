library verilog;
use verilog.vl_types.all;
entity NanoProc_vlg_vec_tst is
end NanoProc_vlg_vec_tst;
