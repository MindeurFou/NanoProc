package pgm_def is
type T_ROMPGM is array (integer range 0 to 99) of integer range 0 to 2**24-1;
constant ROMPGM : T_ROMPGM := (
16#C02400#,16#801000#,16#C0A040#,16#000103#,16#00004C#,16#000018#,16#20495E#,16#C01B03#,
16#AFFD5E#,16#401003#,16#C0020E#,16#C002C0#,16#00030F#,16#8005C0#,16#40050E#,16#00405E#,
16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,
16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,
16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,
16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,
16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,
16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,
16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,
16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,16#00001D#,
16#C04880#,16#C0CCC0#,16#000383#,16#802180#,16#C0149C#,16#2FABDE#,16#C01080#,16#C001C0#,
16#000385#,16#802080#,16#C0028E#,16#C005D4#,16#0002D5#,16#400255#,16#000255#,16#C00255#,
16#00011E#,16#00005E#,16#0FFF5E#,16#0FFE5E#);
end package;

----------------------
-- Source du fichier :
-- ;Exemple de fichier source assembleur NanoCPU
-- 
-- 
--    MOVE W0,#0x24  ; Charge 24H dans W0
-- TOTO: EQU 0x5
-- 
-- DEB:
--    MOVE MEM,W0   ; Range W0 � l'adresse 10h
--    MOVE W1,#0xA0  ; Charge A0H dans W1
--    ADD W0,W1      ; W0<-W0+W1
--    INC W1
--    SETC
--    ;DEC 0x21B  ; ill�gal
-- LBL1: beq lbl2
--    ADD W0,#0x1B   ;
--    BMI LBL1       ;
--    ADD W0,0x10    ;
--    ROL W0,#2
--    MOVE W3,#2
--    ROR W0,W3
--    MOVE 0x05,W3
--    ROL W0,0x05
--    bra lbl2
--    ORG 0x50
-- lbl2:
--    MOVE W2,#0x48
--    MOVE W3,#0b11001100
--    ADD W2,W3
--    MOVE 0x21,W2
--    CMP W2,#0x14
--    BEQ DEB
--    MOVE W2,#0x10
--    MOVE W3,#0x01
--    ADDC W2,W3
--    MOVE 0x20,W2
--    ROL W2,#2
--    BCLR W3,#5
--    BSET W3,W2
--    BSET W1,0x2
--    BSET W1,W2
--    BSET W1,#2
--    JMP DEB        ; {.opbr=BR,.cond=ALWS,.mode=ABS,.dest=1},
--    bra fin
-- fin: bra fin
--    bra fin
-- ;   ADD 0x12,W3    ; interdit !
-- MEM: EQU 0x10
-- 
-- 
