library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ProcTest is
end entity;

architecture behav of ProcTest is
component FemtoProc is
   port(
      clk, raz : in bit;
-- signaux de debug :
      RomData: out std_logic_vector(23 downto 0);
      AdRAM : in std_logic_vector(7 downto 0);
      RamData: out std_logic_vector(7 downto 0);
      NumReg: in std_logic_vector(1 downto 0);
      RegOut: out std_logic_vector(7 downto 0);
      PCOut: out std_logic_vector(11 downto 0);
      Zout,Cout,Nout,Vout: out std_logic
   );
   end component;

signal clk : bit:='0';
signal raz : bit:='1';
signal RomData: std_logic_vector(23 downto 0):=(others=>'0');
signal AdRAM : std_logic_vector(7 downto 0):=(others=>'0');
signal RamData: std_logic_vector(7 downto 0):=(others=>'0');
signal NumReg: std_logic_vector(1 downto 0):=(others=>'0');
signal RegOut: std_logic_vector(7 downto 0):=(others=>'0');
signal PCOut: std_logic_vector(11 downto 0):=(others=>'0');
signal Zout,Cout,Nout,Vout: std_logic;

function v2hex(v:std_logic_vector(3 downto 0)) return string is
constant t : string (1 to 16) := "0123456789ABCDEF";
variable h : string(1 to 1);
variable n : integer range 1 to 16;
begin
   n:=to_integer(unsigned(v))+1;
   return t(n to n);
end function;

function vv2hex(v:std_logic_vector) return string is
variable h:string(1 to v'length/4);
variable n: integer range 0 to v'length;
begin
   for i in 0 to v'length/4-1 loop
   n:=v'length-1-4*i;
   h(i+1 to i+1):=v2hex(v(n downto n-3));
   end loop;
   return h;
end function;

function b2str(b: std_logic) return string is
begin
  if b='0' then return "0";
  else return "1";
  end if;
end function;

begin
   process
   begin
   raz<='1'; wait for 10 ns; raz<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (C02400)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"001" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"24" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (801000)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"002" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"24" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   AdRAM<=X"10";
   wait for 1 ns;
   assert RamData=X"24" report "Erreur (010)<-W0";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (C0A040)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"003" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"24" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A0" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (000103)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"004" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"C4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A0" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":INC (00004C)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"005" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"C4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":SETC (000018)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"006" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"C4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BEQ (20495E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"007" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"C4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (C01B03)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"008" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"DF" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BMI (AFFD5E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"006" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"DF" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BEQ (20495E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"007" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"DF" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (C01B03)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"008" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"FA" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BMI (AFFD5E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"006" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"FA" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BEQ (20495E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"007" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"FA" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (C01B03)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"008" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"15" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BMI (AFFD5E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"009" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"15" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (401003)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"00A" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"39" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ROL (C0020E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"00B" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (C002C0)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"00C" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"02" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ROR (00030F)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"00D" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"39" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"02" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (8005C0)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"00E" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"39" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"02" report "Erreur W3";
   AdRAM<=X"05";
   wait for 1 ns;
   assert RamData=X"02" report "Erreur (005)<-W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ROL (40050E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"00F" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"02" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BRA (00405E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"050" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"00" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"02" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (C04880)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"051" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"48" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"02" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (C0CCC0)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"052" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"48" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (000383)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"053" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (802180)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"054" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   AdRAM<=X"21";
   wait for 1 ns;
   assert RamData=X"14" report "Erreur (021)<-W2";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":CMP (C0149C)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"055" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='1' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BEQ (2FABDE)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"001" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='1' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (801000)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"002" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   AdRAM<=X"10";
   wait for 1 ns;
   assert RamData=X"E4" report "Erreur (010)<-W0";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":MOVE (C0A040)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"003" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"E4" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A0" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (000103)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"004" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"84" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A0" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":INC (00004C)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"005" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"84" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":SETC (000018)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"006" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"84" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BEQ (20495E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"007" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"84" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (C01B03)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"008" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"9F" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BMI (AFFD5E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"006" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"9F" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BEQ (20495E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"007" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"9F" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (C01B03)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"008" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"BA" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BMI (AFFD5E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"006" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"BA" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BEQ (20495E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"007" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"BA" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (C01B03)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"008" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"D5" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BMI (AFFD5E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"006" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"D5" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BEQ (20495E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"007" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"D5" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (C01B03)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"008" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"F0" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BMI (AFFD5E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"006" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"F0" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BEQ (20495E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"007" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"F0" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (C01B03)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"008" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"0B" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":BMI (AFFD5E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"009" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='0' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"0B" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ADD (401003)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"00A" report "Erreur PC";
   assert COut='0' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"EF" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
   report vv2hex(PCOut)&":ROL (C0020E)";
   clk<='1'; wait for 10 ns;
   report "C="&b2str(COut)&" Z="&b2str(ZOut)&" N="&b2str(NOut)&" V="&b2str(VOut);
   assert PCOut=X"00B" report "Erreur PC";
   assert COut='1' report "Erreur C";
   assert ZOut='0' report "Erreur Z";
   assert NOut='1' report "Erreur N";
   assert VOut='0' report "Erreur V";
   NumReg<="00";
   wait for 1 ns;
   assert RegOut=X"BD" report "Erreur W0";
   NumReg<="01";
   wait for 1 ns;
   assert RegOut=X"A1" report "Erreur W1";
   NumReg<="10";
   wait for 1 ns;
   assert RegOut=X"14" report "Erreur W2";
   NumReg<="11";
   wait for 1 ns;
   assert RegOut=X"CC" report "Erreur W3";
   clk<='0'; wait for 10 ns;
wait;
end process;
u1: FemtoProc port map(clk,raz,RomData,AdRAM,RamData,NumReg,RegOut,PCOut,Zout,Cout,Nout,Vout);
end architecture;
